LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY q5 IS
	PORT (a, b, s   : IN SIGNED(3 downto 0);
	      m, ci     : IN STD_LOGIC;
	      f         : OUT SIGNED(3 downto 0);
	      p, g      : OUT STD_LOGIC;
	      aeqb, cn4 : OUT STD_LOGIC);
END q5;

ARCHITECTURE struct OF q5 IS
BEGIN
END struct;
