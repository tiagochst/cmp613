LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.NUMERIC_STD.all;
USE work.PAC_DEFS.all;
  
PACKAGE pac_sprites IS  
  --Desenhos do pacman nas quatro possiveis direcoes
  CONSTANT PAC_BLKMAPS: t_ovl_blk_dir_vet := (
  CIMA =>   ((BLK_PAC_CIM_00, BLK_PAC_CIM_01, BLK_PAC_CIM_02, BLK_PAC_CIM_03, BLK_PAC_CIM_04),
             (BLK_PAC_CIM_10, BLK_PAC_CIM_11, BLK_PAC_CIM_12, BLK_PAC_CIM_13, BLK_PAC_CIM_14),
             (BLK_PAC_CIM_20, BLK_PAC_CIM_21, BLK_PAC_CIM_22, BLK_PAC_CIM_23, BLK_PAC_CIM_24),
             (BLK_PAC_CIM_30, BLK_PAC_CIM_31, BLK_PAC_CIM_32, BLK_PAC_CIM_33, BLK_PAC_CIM_34),
             (BLK_PAC_CIM_40, BLK_PAC_CIM_41, BLK_PAC_CIM_42, BLK_PAC_CIM_43, BLK_PAC_CIM_44)),
  DIREI =>  ((BLK_PAC_DIR_00, BLK_PAC_DIR_01, BLK_PAC_DIR_02, BLK_PAC_DIR_03, BLK_PAC_DIR_04),
             (BLK_PAC_DIR_10, BLK_PAC_DIR_11, BLK_PAC_DIR_12, BLK_PAC_DIR_13, BLK_PAC_DIR_14),
             (BLK_PAC_DIR_20, BLK_PAC_DIR_21, BLK_PAC_DIR_22, BLK_PAC_DIR_23, BLK_PAC_DIR_24),
             (BLK_PAC_DIR_30, BLK_PAC_DIR_31, BLK_PAC_DIR_32, BLK_PAC_DIR_33, BLK_PAC_DIR_34),
             (BLK_PAC_DIR_40, BLK_PAC_DIR_41, BLK_PAC_DIR_42, BLK_PAC_DIR_43, BLK_PAC_DIR_44)),
    BAIXO =>  ((BLK_PAC_BAI_00, BLK_PAC_BAI_01, BLK_PAC_BAI_02, BLK_PAC_BAI_03, BLK_PAC_BAI_04),
             (BLK_PAC_BAI_10, BLK_PAC_BAI_11, BLK_PAC_BAI_12, BLK_PAC_BAI_13, BLK_PAC_BAI_14),
             (BLK_PAC_BAI_20, BLK_PAC_BAI_21, BLK_PAC_BAI_22, BLK_PAC_BAI_23, BLK_PAC_BAI_24),
             (BLK_PAC_BAI_30, BLK_PAC_BAI_31, BLK_PAC_BAI_32, BLK_PAC_BAI_33, BLK_PAC_BAI_34),
             (BLK_PAC_BAI_40, BLK_PAC_BAI_41, BLK_PAC_BAI_42, BLK_PAC_BAI_43, BLK_PAC_BAI_44)),
  ESQUE =>  ((BLK_PAC_ESQ_00, BLK_PAC_ESQ_01, BLK_PAC_ESQ_02, BLK_PAC_ESQ_03, BLK_PAC_ESQ_04),
             (BLK_PAC_ESQ_10, BLK_PAC_ESQ_11, BLK_PAC_ESQ_12, BLK_PAC_ESQ_13, BLK_PAC_ESQ_14),
             (BLK_PAC_ESQ_20, BLK_PAC_ESQ_21, BLK_PAC_ESQ_22, BLK_PAC_ESQ_23, BLK_PAC_ESQ_24),
             (BLK_PAC_ESQ_30, BLK_PAC_ESQ_31, BLK_PAC_ESQ_32, BLK_PAC_ESQ_33, BLK_PAC_ESQ_34),
             (BLK_PAC_ESQ_40, BLK_PAC_ESQ_41, BLK_PAC_ESQ_42, BLK_PAC_ESQ_43, BLK_PAC_ESQ_44)),
  OTHERS => (OTHERS => (OTHERS => BLK_NULL))
  );
  
  CONSTANT PAC_FECH_BLKMAP: t_ovl_blk_5x5 := (
    (BLK_PAC_FECH_00, BLK_PAC_FECH_01, BLK_PAC_FECH_02, BLK_PAC_FECH_03, BLK_PAC_FECH_04),
    (BLK_PAC_FECH_10, BLK_PAC_FECH_11, BLK_PAC_FECH_12, BLK_PAC_FECH_13, BLK_PAC_FECH_14),
    (BLK_PAC_FECH_20, BLK_PAC_FECH_21, BLK_PAC_FECH_22, BLK_PAC_FECH_23, BLK_PAC_FECH_24),
    (BLK_PAC_FECH_30, BLK_PAC_FECH_31, BLK_PAC_FECH_32, BLK_PAC_FECH_33, BLK_PAC_FECH_34),
    (BLK_PAC_FECH_40, BLK_PAC_FECH_41, BLK_PAC_FECH_42, BLK_PAC_FECH_43, BLK_PAC_FECH_44));

  CONSTANT PAC_FECV_BLKMAP: t_ovl_blk_5x5 := (
    (BLK_PAC_FECV_00, BLK_PAC_FECV_01, BLK_PAC_FECV_02, BLK_PAC_FECV_03, BLK_PAC_FECV_04),
    (BLK_PAC_FECV_10, BLK_PAC_FECV_11, BLK_PAC_FECV_12, BLK_PAC_FECV_13, BLK_PAC_FECV_14),
    (BLK_PAC_FECV_20, BLK_PAC_FECV_21, BLK_PAC_FECV_22, BLK_PAC_FECV_23, BLK_PAC_FECV_24),
    (BLK_PAC_FECV_30, BLK_PAC_FECV_31, BLK_PAC_FECV_32, BLK_PAC_FECV_33, BLK_PAC_FECV_34),
    (BLK_PAC_FECV_40, BLK_PAC_FECV_41, BLK_PAC_FECV_42, BLK_PAC_FECV_43, BLK_PAC_FECV_44));
    
  CONSTANT FAN_BLKMAPS: t_fans_ovl_blk_dir_vet := (
  0 => ( --primeiro fantasma:
  CIMA =>  ((BLK_FAN_GRN_00,     BLK_FAN_GRN_01,     BLK_FAN_GRN_02,     BLK_FAN_GRN_03, BLK_FAN_GRN_04),
       (BLK_FAN_GRN_10, BLK_EYE_GRN_CIM_00, BLK_EYE_GRN_CIM_01, BLK_EYE_GRN_CIM_02, BLK_FAN_GRN_14),
       (BLK_FAN_GRN_20, BLK_EYE_GRN_CIM_10, BLK_EYE_GRN_CIM_11, BLK_EYE_GRN_CIM_12, BLK_FAN_GRN_24),
       (BLK_FAN_GRN_30,     BLK_FAN_GRN_31,     BLK_FAN_GRN_32,     BLK_FAN_GRN_33, BLK_FAN_GRN_34),
       (BLK_FAN_GRN_40,     BLK_FAN_GRN_41,     BLK_FAN_GRN_42,     BLK_FAN_GRN_43, BLK_FAN_GRN_44)),
  DIREI=> ((BLK_FAN_GRN_00,     BLK_FAN_GRN_01,     BLK_FAN_GRN_02,     BLK_FAN_GRN_03, BLK_FAN_GRN_04),
       (BLK_FAN_GRN_10, BLK_EYE_GRN_DIR_00, BLK_EYE_GRN_DIR_01, BLK_EYE_GRN_DIR_02, BLK_FAN_GRN_14),
       (BLK_FAN_GRN_20, BLK_EYE_GRN_DIR_10, BLK_EYE_GRN_DIR_11, BLK_EYE_GRN_DIR_12, BLK_FAN_GRN_24),
       (BLK_FAN_GRN_30,     BLK_FAN_GRN_31,     BLK_FAN_GRN_32,     BLK_FAN_GRN_33, BLK_FAN_GRN_34),
       (BLK_FAN_GRN_40,     BLK_FAN_GRN_41,     BLK_FAN_GRN_42,     BLK_FAN_GRN_43, BLK_FAN_GRN_44)),
  BAIXO=>  ((BLK_FAN_GRN_00,     BLK_FAN_GRN_01,     BLK_FAN_GRN_02,     BLK_FAN_GRN_03, BLK_FAN_GRN_04),
       (BLK_FAN_GRN_10, BLK_EYE_GRN_BAI_00, BLK_EYE_GRN_BAI_01, BLK_EYE_GRN_BAI_02, BLK_FAN_GRN_14),
       (BLK_FAN_GRN_20, BLK_EYE_GRN_BAI_10, BLK_EYE_GRN_BAI_11, BLK_EYE_GRN_BAI_12, BLK_FAN_GRN_24),
       (BLK_FAN_GRN_30,     BLK_FAN_GRN_31,     BLK_FAN_GRN_32,     BLK_FAN_GRN_33, BLK_FAN_GRN_34),
       (BLK_FAN_GRN_40,     BLK_FAN_GRN_41,     BLK_FAN_GRN_42,     BLK_FAN_GRN_43, BLK_FAN_GRN_44)),
  ESQUE=>  ((BLK_FAN_GRN_00,     BLK_FAN_GRN_01,     BLK_FAN_GRN_02,     BLK_FAN_GRN_03, BLK_FAN_GRN_04),
       (BLK_FAN_GRN_10, BLK_EYE_GRN_ESQ_00, BLK_EYE_GRN_ESQ_01, BLK_EYE_GRN_ESQ_02, BLK_FAN_GRN_14),
       (BLK_FAN_GRN_20, BLK_EYE_GRN_ESQ_10, BLK_EYE_GRN_ESQ_11, BLK_EYE_GRN_ESQ_12, BLK_FAN_GRN_24),
       (BLK_FAN_GRN_30,     BLK_FAN_GRN_31,     BLK_FAN_GRN_32,     BLK_FAN_GRN_33, BLK_FAN_GRN_34),
       (BLK_FAN_GRN_40,     BLK_FAN_GRN_41,     BLK_FAN_GRN_42,     BLK_FAN_GRN_43, BLK_FAN_GRN_44)),
  OTHERS => (OTHERS => (OTHERS => BLK_NULL))),
  1 => ( --segundo fantasma:
  CIMA =>  ((BLK_FAN_RED_00,     BLK_FAN_RED_01,     BLK_FAN_RED_02,     BLK_FAN_RED_03, BLK_FAN_RED_04),
       (BLK_FAN_RED_10, BLK_EYE_RED_CIM_00, BLK_EYE_RED_CIM_01, BLK_EYE_RED_CIM_02, BLK_FAN_RED_14),
       (BLK_FAN_RED_20, BLK_EYE_RED_CIM_10, BLK_EYE_RED_CIM_11, BLK_EYE_RED_CIM_12, BLK_FAN_RED_24),
       (BLK_FAN_RED_30,     BLK_FAN_RED_31,     BLK_FAN_RED_32,     BLK_FAN_RED_33, BLK_FAN_RED_34),
       (BLK_FAN_RED_40,     BLK_FAN_RED_41,     BLK_FAN_RED_42,     BLK_FAN_RED_43, BLK_FAN_RED_44)),
  DIREI=> ((BLK_FAN_RED_00,     BLK_FAN_RED_01,     BLK_FAN_RED_02,     BLK_FAN_RED_03, BLK_FAN_RED_04),
       (BLK_FAN_RED_10, BLK_EYE_RED_DIR_00, BLK_EYE_RED_DIR_01, BLK_EYE_RED_DIR_02, BLK_FAN_RED_14),
       (BLK_FAN_RED_20, BLK_EYE_RED_DIR_10, BLK_EYE_RED_DIR_11, BLK_EYE_RED_DIR_12, BLK_FAN_RED_24),
       (BLK_FAN_RED_30,     BLK_FAN_RED_31,     BLK_FAN_RED_32,     BLK_FAN_RED_33, BLK_FAN_RED_34),
       (BLK_FAN_RED_40,     BLK_FAN_RED_41,     BLK_FAN_RED_42,     BLK_FAN_RED_43, BLK_FAN_RED_44)),
  BAIXO=>  ((BLK_FAN_RED_00,     BLK_FAN_RED_01,     BLK_FAN_RED_02,     BLK_FAN_RED_03, BLK_FAN_RED_04),
       (BLK_FAN_RED_10, BLK_EYE_RED_BAI_00, BLK_EYE_RED_BAI_01, BLK_EYE_RED_BAI_02, BLK_FAN_RED_14),
       (BLK_FAN_RED_20, BLK_EYE_RED_BAI_10, BLK_EYE_RED_BAI_11, BLK_EYE_RED_BAI_12, BLK_FAN_RED_24),
       (BLK_FAN_RED_30,     BLK_FAN_RED_31,     BLK_FAN_RED_32,     BLK_FAN_RED_33, BLK_FAN_RED_34),
       (BLK_FAN_RED_40,     BLK_FAN_RED_41,     BLK_FAN_RED_42,     BLK_FAN_RED_43, BLK_FAN_RED_44)),
  ESQUE=>  ((BLK_FAN_RED_00,     BLK_FAN_RED_01,     BLK_FAN_RED_02,     BLK_FAN_RED_03, BLK_FAN_RED_04),
       (BLK_FAN_RED_10, BLK_EYE_RED_ESQ_00, BLK_EYE_RED_ESQ_01, BLK_EYE_RED_ESQ_02, BLK_FAN_RED_14),
       (BLK_FAN_RED_20, BLK_EYE_RED_ESQ_10, BLK_EYE_RED_ESQ_11, BLK_EYE_RED_ESQ_12, BLK_FAN_RED_24),
       (BLK_FAN_RED_30,     BLK_FAN_RED_31,     BLK_FAN_RED_32,     BLK_FAN_RED_33, BLK_FAN_RED_34),
       (BLK_FAN_RED_40,     BLK_FAN_RED_41,     BLK_FAN_RED_42,     BLK_FAN_RED_43, BLK_FAN_RED_44)),
  OTHERS => (OTHERS => (OTHERS => BLK_NULL)))
  );
  
  CONSTANT FAN_DEAD_BLKMAPS: t_ovl_blk_dir_vet := (
  CIMA =>  ((  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_CIM_00, BLK_EYE_BLK_CIM_01, BLK_EYE_BLK_CIM_02,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_CIM_10, BLK_EYE_BLK_CIM_11, BLK_EYE_BLK_CIM_12,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL)),
  DIREI=> ((  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_DIR_00, BLK_EYE_BLK_DIR_01, BLK_EYE_BLK_DIR_02,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_DIR_10, BLK_EYE_BLK_DIR_11, BLK_EYE_BLK_DIR_12,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL)),
  BAIXO=>  ((  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_BAI_00, BLK_EYE_BLK_BAI_01, BLK_EYE_BLK_BAI_02,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_BAI_10, BLK_EYE_BLK_BAI_11, BLK_EYE_BLK_BAI_12,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL)),
  ESQUE=>  ((  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_ESQ_00, BLK_EYE_BLK_ESQ_01, BLK_EYE_BLK_ESQ_02,   BLK_NULL),
       (  BLK_NULL, BLK_EYE_BLK_ESQ_10, BLK_EYE_BLK_ESQ_11, BLK_EYE_BLK_ESQ_12,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL),
       (  BLK_NULL,       BLK_NULL,       BLK_NULL,       BLK_NULL,   BLK_NULL)),
  OTHERS => (OTHERS => (OTHERS => BLK_NULL))
  );
  
  CONSTANT FAN_VULN_BLKMAP: t_ovl_blk_5x5 := (
    (BLK_FAN_VULN_00, BLK_FAN_VULN_01, BLK_FAN_VULN_02, BLK_FAN_VULN_03, BLK_FAN_VULN_04),
    (BLK_FAN_VULN_10, BLK_FAN_VULN_11, BLK_FAN_VULN_12, BLK_FAN_VULN_13, BLK_FAN_VULN_14),
    (BLK_FAN_VULN_20, BLK_FAN_VULN_21, BLK_FAN_VULN_22, BLK_FAN_VULN_23, BLK_FAN_VULN_24),
    (BLK_FAN_VULN_30, BLK_FAN_VULN_31, BLK_FAN_VULN_32, BLK_FAN_VULN_33, BLK_FAN_VULN_34),
    (BLK_FAN_VULN_40, BLK_FAN_VULN_41, BLK_FAN_VULN_42, BLK_FAN_VULN_43, BLK_FAN_VULN_44));
    
  CONSTANT FRUTA_BLKMAP: t_frut_ovl_blk_vet := (
    1 =>((BLK_MACA_00, BLK_MACA_01, BLK_MACA_02, BLK_MACA_03, BLK_MACA_04),
      (BLK_MACA_10, BLK_MACA_11, BLK_MACA_12, BLK_MACA_13, BLK_MACA_14),
      (BLK_MACA_20, BLK_MACA_21, BLK_MACA_22, BLK_MACA_23, BLK_MACA_24),
      (BLK_MACA_30, BLK_MACA_31, BLK_MACA_32, BLK_MACA_33, BLK_MACA_34),
      (BLK_MACA_40, BLK_MACA_41, BLK_MACA_42, BLK_MACA_43, BLK_MACA_44)),
    2 =>((BLK_CEREJA_00, BLK_CEREJA_01, BLK_CEREJA_02, BLK_CEREJA_03, BLK_CEREJA_04),
      (BLK_CEREJA_10, BLK_CEREJA_11, BLK_CEREJA_12, BLK_CEREJA_13, BLK_CEREJA_14),
      (BLK_CEREJA_20, BLK_CEREJA_21, BLK_CEREJA_22, BLK_CEREJA_23, BLK_CEREJA_24),
      (BLK_CEREJA_30, BLK_CEREJA_31, BLK_CEREJA_32, BLK_CEREJA_33, BLK_CEREJA_34),
      (BLK_CEREJA_40, BLK_CEREJA_41, BLK_CEREJA_42, BLK_CEREJA_43, BLK_CEREJA_44)),
    OTHERS => (OTHERS => (OTHERS => BLK_NULL))
  );
  
  CONSTANT SPRITES_RED: t_sprite5_vet := (
  BLK_COIN       => ("00000","01110","01110","01110","00000"),
  BLK_SPC_COIN    => ("11111","11111","11111","11111","11111"),  
  BLK_DOOR    => ("11111","11111","11111","00000","00000"),
  OTHERS      => (OTHERS => (OTHERS => '0')));
  
  CONSTANT SPRITES_GRN: t_sprite5_vet := (
  BLK_COIN      => ("00000","01110","01110","01110","00000"),
  BLK_SPC_COIN    => ("11111","11111","11111","11111","11111"),
  OTHERS      => (OTHERS => (OTHERS => '0')));
  
  CONSTANT SPRITES_BLU: t_sprite5_vet := (
  BLK_COIN       => ("00000","01110","01110","01110","00000"),
  BLK_SPC_COIN    => ("11111","11111","11111","11111","11111"),
  BLK_WALL_V     => ("10010","10010","10010","10010","10010"),
  BLK_WALL_H     => ("11111","00000","00000","11111","00000"),
  BLK_WALL_Q      => ("00111","01100","11000","10001","10010"),
  BLK_WALL_W      => ("11000","01100","00110","00010","10010"),
  BLK_WALL_E      => ("10001","11000","01100","00111","00000"),
  BLK_WALL_R      => ("00010","00110","01100","11000","00000"),
  OTHERS      => (OTHERS => (OTHERS => '0')));

  CONSTANT OVL_SPRITES_RED: t_ovl_sprite5_vet := (
  BLK_PAC_CIM_00 => ("00000","00000","00000","00000","00001"),
  BLK_PAC_CIM_01 => ("00000","00000","00000","11000","11000"),
  BLK_PAC_CIM_02 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_03 => ("00000","00000","00000","00011","00011"),
  BLK_PAC_CIM_04 => ("00000","00000","00000","00000","10000"),
  BLK_PAC_CIM_10 => ("00011","00111","00111","01111","01111"),
  BLK_PAC_CIM_11 => ("11100","11100","11110","11110","11111"),
  BLK_PAC_CIM_12 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_13 => ("00111","00111","01111","01111","11111"),
  BLK_PAC_CIM_14 => ("11000","11100","11100","11110","11110"),
  BLK_PAC_CIM_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_CIM_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_22 => ("10001","10001","11011","11111","11111"),
  BLK_PAC_CIM_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_CIM_30 => ("00111","00111","00011","00001","00000"),
  BLK_PAC_CIM_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_34 => ("11100","11100","11000","10000","00000"),
  BLK_PAC_CIM_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_41 => ("01111","00011","00001","00000","00000"),
  BLK_PAC_CIM_42 => ("11111","11111","11111","00000","00000"),
  BLK_PAC_CIM_43 => ("11110","11000","10000","00000","00000"),
  BLK_PAC_CIM_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_01 => ("00000","00000","00011","00111","01111"),
  BLK_PAC_DIR_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_DIR_03 => ("00000","11000","11110","11111","11111"),
  BLK_PAC_DIR_04 => ("00000","00000","00000","00000","10000"),
  BLK_PAC_DIR_10 => ("00000","00001","00001","00011","00111"),
  BLK_PAC_DIR_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_13 => ("11111","11111","11111","11100","10000"),
  BLK_PAC_DIR_14 => ("11000","11000","00000","00000","00000"),
  BLK_PAC_DIR_20 => ("00111","00111","00111","00111","00111"),
  BLK_PAC_DIR_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_22 => ("11111","11100","11000","11100","11111"),
  BLK_PAC_DIR_23 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_24 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_30 => ("00111","00011","00001","00001","00000"),
  BLK_PAC_DIR_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_33 => ("10000","11100","11111","11111","11111"),
  BLK_PAC_DIR_34 => ("00000","00000","00000","11000","11000"),
  BLK_PAC_DIR_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_41 => ("01111","00111","00011","00000","00000"),
  BLK_PAC_DIR_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_DIR_43 => ("11111","11111","11110","11000","00000"),
  BLK_PAC_DIR_44 => ("10000","00000","00000","00000","00000"),
  BLK_PAC_BAI_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_01 => ("00000","00000","00001","00011","01111"),
  BLK_PAC_BAI_02 => ("00000","00000","11111","11111","11111"),
  BLK_PAC_BAI_03 => ("00000","00000","10000","11000","11110"),
  BLK_PAC_BAI_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_10 => ("00000","00001","00011","00111","00111"),
  BLK_PAC_BAI_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_14 => ("00000","10000","11000","11100","11100"),
  BLK_PAC_BAI_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_BAI_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_22 => ("11111","11111","11011","10001","10001"),
  BLK_PAC_BAI_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_BAI_30 => ("01111","01111","00111","00111","00011"),
  BLK_PAC_BAI_31 => ("11111","11110","11110","11100","11100"),
  BLK_PAC_BAI_32 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_33 => ("11111","01111","01111","00111","00111"),
  BLK_PAC_BAI_34 => ("11110","11110","11100","11100","11000"),
  BLK_PAC_BAI_40 => ("00001","00000","00000","00000","00000"),
  BLK_PAC_BAI_41 => ("11000","11000","00000","00000","00000"),
  BLK_PAC_BAI_42 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_43 => ("00011","00011","00000","00000","00000"),
  BLK_PAC_BAI_44 => ("10000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_00 => ("00000","00000","00000","00000","00001"),
  BLK_PAC_ESQ_01 => ("00000","00011","01111","11111","11111"),
  BLK_PAC_ESQ_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_ESQ_03 => ("00000","00000","11000","11100","11110"),
  BLK_PAC_ESQ_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_10 => ("00011","00011","00000","00000","00000"),
  BLK_PAC_ESQ_11 => ("11111","11111","11111","00111","00001"),
  BLK_PAC_ESQ_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_14 => ("00000","10000","10000","11000","11100"),
  BLK_PAC_ESQ_20 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_21 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_22 => ("11111","00111","00011","00111","11111"),
  BLK_PAC_ESQ_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_24 => ("11100","11100","11100","11100","11100"),
  BLK_PAC_ESQ_30 => ("00000","00000","00000","00011","00011"),
  BLK_PAC_ESQ_31 => ("00001","00111","11111","11111","11111"),
  BLK_PAC_ESQ_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_34 => ("11100","11000","10000","10000","00000"),
  BLK_PAC_ESQ_40 => ("00001","00000","00000","00000","00000"),
  BLK_PAC_ESQ_41 => ("11111","11111","01111","00011","00000"),
  BLK_PAC_ESQ_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_ESQ_43 => ("11110","11100","11000","00000","00000"),
  BLK_PAC_ESQ_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_01 => ("00000","00000","00001","00011","01111"),
  BLK_PAC_FECV_02 => ("00000","00000","11111","11111","11111"),
  BLK_PAC_FECV_03 => ("00000","00000","10000","11000","11110"),
  BLK_PAC_FECV_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_10 => ("00000","00001","00011","00111","00111"),
  BLK_PAC_FECV_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_14 => ("00000","10000","11000","11100","11100"),
  BLK_PAC_FECV_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_FECV_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_22 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_FECV_30 => ("00111","00111","00011","00001","00000"),
  BLK_PAC_FECV_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_34 => ("11100","11100","11000","10000","00000"),
  BLK_PAC_FECV_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_41 => ("01111","00011","00001","00000","00000"),
  BLK_PAC_FECV_42 => ("11111","11111","11111","00000","00000"),
  BLK_PAC_FECV_43 => ("11110","11000","10000","00000","00000"),
  BLK_PAC_FECV_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_01 => ("00000","00000","00011","00111","01111"),
  BLK_PAC_FECH_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_FECH_03 => ("00000","00000","11000","11100","11110"),
  BLK_PAC_FECH_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_10 => ("00000","00001","00001","00011","00111"),
  BLK_PAC_FECH_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_14 => ("00000","10000","10000","11000","11100"),
  BLK_PAC_FECH_20 => ("00111","00111","00111","00111","00111"),
  BLK_PAC_FECH_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_22 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_24 => ("11100","11100","11100","11100","11100"),
  BLK_PAC_FECH_30 => ("00111","00011","00001","00001","00000"),
  BLK_PAC_FECH_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_34 => ("11100","11000","10000","10000","00000"),
  BLK_PAC_FECH_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_41 => ("01111","00111","00011","00000","00000"),
  BLK_PAC_FECH_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_FECH_43 => ("11110","11100","11000","00000","00000"),
  BLK_PAC_FECH_44 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_RED_00 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_RED_01 => ("00000","00111","01111","11111","11111"),
  BLK_FAN_RED_02 => ("00000","11111","11111","11111","11111"),
  BLK_FAN_RED_03 => ("00000","11000","11100","11110","11110"),
  BLK_FAN_RED_04 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_RED_10 => ("00001","00011","00011","00111","00111"),
  BLK_FAN_RED_14 => ("00000","10000","10000","11000","11000"),
  BLK_FAN_RED_20 => ("00111","00111","01111","01111","01111"),
  BLK_FAN_RED_24 => ("11000","11000","11100","11100","11100"),
  BLK_FAN_RED_30 => ("01111","01111","01111","01111","01111"),
  BLK_FAN_RED_31 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_RED_32 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_RED_33 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_RED_34 => ("11100","11100","11100","11100","11100"),
  BLK_FAN_RED_40 => ("01111","01111","01111","00110","00000"),
  BLK_FAN_RED_41 => ("10011","00001","00000","00000","00000"),
  BLK_FAN_RED_42 => ("11111","11111","11110","01100","00000"),
  BLK_FAN_RED_43 => ("10011","00001","00001","00000","00000"),
  BLK_FAN_RED_44 => ("11100","11100","11100","11000","00000"),
  BLK_EYE_RED_CIM_00 => ("10001","10001","10001","11111","11111"),
  BLK_EYE_RED_CIM_01 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_CIM_02 => ("00011","00011","00011","11111","11111"),
  BLK_EYE_RED_CIM_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_CIM_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_CIM_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_DIR_00 => ("11111","11111","11100","11100","11100"),
  BLK_EYE_RED_DIR_01 => ("11111","11111","01111","01111","01111"),
  BLK_EYE_RED_DIR_02 => ("11111","11111","11000","11000","11000"),
  BLK_EYE_RED_DIR_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_DIR_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_DIR_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_BAI_00 => ("11111","11111","11111","11111","11000"),
  BLK_EYE_RED_BAI_01 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_BAI_02 => ("11111","11111","11111","11111","10001"),
  BLK_EYE_RED_BAI_10 => ("11000","11000","11111","11111","11111"),
  BLK_EYE_RED_BAI_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_BAI_12 => ("10001","10001","11111","11111","11111"),
  BLK_EYE_RED_ESQ_00 => ("11111","11111","00011","00011","00011"),
  BLK_EYE_RED_ESQ_01 => ("11111","11111","11110","11110","11110"),
  BLK_EYE_RED_ESQ_02 => ("11111","11111","00111","00111","00111"),
  BLK_EYE_RED_ESQ_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_ESQ_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_RED_ESQ_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_00 => ("00001","10001","10001","11111","11111"),
  BLK_EYE_GRN_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_CIM_02 => ("00010","00011","00011","11111","11111"),
  BLK_EYE_GRN_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_GRN_DIR_00 => ("01111","11111","11100","11100","11100"),
  BLK_EYE_GRN_DIR_01 => ("00000","10001","00001","00001","00001"),
  BLK_EYE_GRN_DIR_02 => ("11110","11111","11000","11000","11000"),
  BLK_EYE_GRN_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_GRN_BAI_00 => ("01111","11111","11111","11111","11000"),
  BLK_EYE_GRN_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_BAI_02 => ("11110","11111","11111","11111","10001"),
  BLK_EYE_GRN_BAI_10 => ("11000","01000","00000","00000","00000"),
  BLK_EYE_GRN_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_BAI_12 => ("10001","10000","00000","00000","00000"),
  BLK_EYE_GRN_ESQ_00 => ("01111","11111","00011","00011","00011"),
  BLK_EYE_GRN_ESQ_01 => ("00000","10001","10000","10000","10000"),
  BLK_EYE_GRN_ESQ_02 => ("11110","11111","00111","00111","00111"),
  BLK_EYE_GRN_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_CIM_00 => ("00001","10001","10001","11111","11111"),
  BLK_EYE_BLK_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_CIM_02 => ("00010","00011","00011","11111","11111"),
  BLK_EYE_BLK_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_DIR_00 => ("01111","11111","11100","11100","11100"),
  BLK_EYE_BLK_DIR_01 => ("00000","10001","00001","00001","00001"),
  BLK_EYE_BLK_DIR_02 => ("11110","11111","11000","11000","11000"),
  BLK_EYE_BLK_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_BAI_00 => ("01111","11111","11111","11111","11000"),
  BLK_EYE_BLK_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_BAI_02 => ("11110","11111","11111","11111","10001"),
  BLK_EYE_BLK_BAI_10 => ("11000","01000","00000","00000","00000"),
  BLK_EYE_BLK_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_BAI_12 => ("10001","10000","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_00 => ("01111","11111","00011","00011","00011"),
  BLK_EYE_BLK_ESQ_01 => ("00000","10001","10000","10000","10000"),
  BLK_EYE_BLK_ESQ_02 => ("11110","11111","00111","00111","00111"),
  BLK_EYE_BLK_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_FAN_VULN_00 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_01 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_02 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_03 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_04 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_10 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_11 => ("00000","00000","00000","00111","00111"),
  BLK_FAN_VULN_12 => ("00000","00000","00000","00001","00001"),
  BLK_FAN_VULN_13 => ("00000","00000","00000","11000","11000"),
  BLK_FAN_VULN_14 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_20 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_21 => ("00111","00000","00000","00000","00000"),
  BLK_FAN_VULN_22 => ("00001","00000","00000","00000","00000"),
  BLK_FAN_VULN_23 => ("11000","00000","00000","00000","00000"),
  BLK_FAN_VULN_24 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_30 => ("00000","00000","00011","00011","00000"),
  BLK_FAN_VULN_31 => ("11100","11100","00011","00011","00000"),
  BLK_FAN_VULN_32 => ("11110","11110","10011","10011","00000"),
  BLK_FAN_VULN_33 => ("01110","01110","10001","10001","00000"),
  BLK_FAN_VULN_34 => ("00000","00000","10000","10000","00000"),
  BLK_FAN_VULN_40 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_41 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_42 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_43 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_44 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_00 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_01 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_02 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_03 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_04 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_10 => ("00000","00000","00000","00001","00011"),
  BLK_MACA_11 => ("00111","01111","11111","11111","11111"),
  BLK_MACA_12 => ("10001","11111","11111","11111","11111"),
  BLK_MACA_13 => ("11100","11110","11111","11111","11111"),
  BLK_MACA_14 => ("00000","00000","00000","10000","11000"),
  BLK_MACA_20 => ("00111","00111","00111","00111","00111"),
  BLK_MACA_21 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_22 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_23 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_24 => ("11100","11100","11100","11100","11100"),
  BLK_MACA_30 => ("00111","00011","00011","00001","00000"),
  BLK_MACA_31 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_32 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_33 => ("11111","11111","11111","11111","11111"),
  BLK_MACA_34 => ("11100","11000","11000","10000","00000"),
  BLK_MACA_40 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_41 => ("01111","00111","00011","00001","00000"),
  BLK_MACA_42 => ("11111","11111","11111","11011","00000"),
  BLK_MACA_43 => ("11110","11100","11000","10000","00000"),
  BLK_MACA_44 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_00 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_01 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_02 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_03 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_04 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_10 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_11 => ("00000","00000","00000","00000","01110"),
  BLK_CEREJA_12 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_13 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_14 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_20 => ("00001","00011","00011","00111","00111"),
  BLK_CEREJA_21 => ("11101","11111","11111","11111","11111"),
  BLK_CEREJA_22 => ("10000","11100","11000","11011","10111"),
  BLK_CEREJA_23 => ("00000","00000","10100","11111","11111"),
  BLK_CEREJA_24 => ("00000","00000","00000","00000","10000"),
  BLK_CEREJA_30 => ("00111","00011","00011","00001","00000"),
  BLK_CEREJA_31 => ("11110","11110","11110","11110","01110"),
  BLK_CEREJA_32 => ("00111","01111","01111","01111","00111"),
  BLK_CEREJA_33 => ("11111","11111","11111","11111","11111"),
  BLK_CEREJA_34 => ("10000","11000","11000","11000","10000"),
  BLK_CEREJA_40 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_41 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_42 => ("00111","00011","00000","00000","00000"),
  BLK_CEREJA_43 => ("11111","11111","11100","00000","00000"),
  BLK_CEREJA_44 => ("10000","00000","00000","00000","00000"),
  OTHERS      => (OTHERS => (OTHERS => '0')));
  
  CONSTANT OVL_SPRITES_GRN: t_ovl_sprite5_vet := (
  BLK_PAC_CIM_00 => ("00000","00000","00000","00000","00001"),
  BLK_PAC_CIM_01 => ("00000","00000","00000","11000","11000"),
  BLK_PAC_CIM_02 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_03 => ("00000","00000","00000","00011","00011"),
  BLK_PAC_CIM_04 => ("00000","00000","00000","00000","10000"),
  BLK_PAC_CIM_10 => ("00011","00111","00111","01111","01111"),
  BLK_PAC_CIM_11 => ("11100","11100","11110","11110","11111"),
  BLK_PAC_CIM_12 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_13 => ("00111","00111","01111","01111","11111"),
  BLK_PAC_CIM_14 => ("11000","11100","11100","11110","11110"),
  BLK_PAC_CIM_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_CIM_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_22 => ("10001","10001","11011","11111","11111"),
  BLK_PAC_CIM_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_CIM_30 => ("00111","00111","00011","00001","00000"),
  BLK_PAC_CIM_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_CIM_34 => ("11100","11100","11000","10000","00000"),
  BLK_PAC_CIM_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_CIM_41 => ("01111","00011","00001","00000","00000"),
  BLK_PAC_CIM_42 => ("11111","11111","11111","00000","00000"),
  BLK_PAC_CIM_43 => ("11110","11000","10000","00000","00000"),
  BLK_PAC_CIM_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_01 => ("00000","00000","00011","00111","01111"),
  BLK_PAC_DIR_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_DIR_03 => ("00000","11000","11110","11111","11111"),
  BLK_PAC_DIR_04 => ("00000","00000","00000","00000","10000"),
  BLK_PAC_DIR_10 => ("00000","00001","00001","00011","00111"),
  BLK_PAC_DIR_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_13 => ("11111","11111","11111","11100","10000"),
  BLK_PAC_DIR_14 => ("11000","11000","00000","00000","00000"),
  BLK_PAC_DIR_20 => ("00111","00111","00111","00111","00111"),
  BLK_PAC_DIR_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_22 => ("11111","11100","11000","11100","11111"),
  BLK_PAC_DIR_23 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_24 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_30 => ("00111","00011","00001","00001","00000"),
  BLK_PAC_DIR_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_DIR_33 => ("10000","11100","11111","11111","11111"),
  BLK_PAC_DIR_34 => ("00000","00000","00000","11000","11000"),
  BLK_PAC_DIR_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_DIR_41 => ("01111","00111","00011","00000","00000"),
  BLK_PAC_DIR_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_DIR_43 => ("11111","11111","11110","11000","00000"),
  BLK_PAC_DIR_44 => ("10000","00000","00000","00000","00000"),
  BLK_PAC_BAI_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_01 => ("00000","00000","00001","00011","01111"),
  BLK_PAC_BAI_02 => ("00000","00000","11111","11111","11111"),
  BLK_PAC_BAI_03 => ("00000","00000","10000","11000","11110"),
  BLK_PAC_BAI_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_10 => ("00000","00001","00011","00111","00111"),
  BLK_PAC_BAI_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_14 => ("00000","10000","11000","11100","11100"),
  BLK_PAC_BAI_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_BAI_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_22 => ("11111","11111","11011","10001","10001"),
  BLK_PAC_BAI_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_BAI_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_BAI_30 => ("01111","01111","00111","00111","00011"),
  BLK_PAC_BAI_31 => ("11111","11110","11110","11100","11100"),
  BLK_PAC_BAI_32 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_33 => ("11111","01111","01111","00111","00111"),
  BLK_PAC_BAI_34 => ("11110","11110","11100","11100","11000"),
  BLK_PAC_BAI_40 => ("00001","00000","00000","00000","00000"),
  BLK_PAC_BAI_41 => ("11000","11000","00000","00000","00000"),
  BLK_PAC_BAI_42 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_BAI_43 => ("00011","00011","00000","00000","00000"),
  BLK_PAC_BAI_44 => ("10000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_00 => ("00000","00000","00000","00000","00001"),
  BLK_PAC_ESQ_01 => ("00000","00011","01111","11111","11111"),
  BLK_PAC_ESQ_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_ESQ_03 => ("00000","00000","11000","11100","11110"),
  BLK_PAC_ESQ_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_10 => ("00011","00011","00000","00000","00000"),
  BLK_PAC_ESQ_11 => ("11111","11111","11111","00111","00001"),
  BLK_PAC_ESQ_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_14 => ("00000","10000","10000","11000","11100"),
  BLK_PAC_ESQ_20 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_21 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_ESQ_22 => ("11111","00111","00011","00111","11111"),
  BLK_PAC_ESQ_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_24 => ("11100","11100","11100","11100","11100"),
  BLK_PAC_ESQ_30 => ("00000","00000","00000","00011","00011"),
  BLK_PAC_ESQ_31 => ("00001","00111","11111","11111","11111"),
  BLK_PAC_ESQ_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_ESQ_34 => ("11100","11000","10000","10000","00000"),
  BLK_PAC_ESQ_40 => ("00001","00000","00000","00000","00000"),
  BLK_PAC_ESQ_41 => ("11111","11111","01111","00011","00000"),
  BLK_PAC_ESQ_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_ESQ_43 => ("11110","11100","11000","00000","00000"),
  BLK_PAC_ESQ_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_01 => ("00000","00000","00001","00011","01111"),
  BLK_PAC_FECV_02 => ("00000","00000","11111","11111","11111"),
  BLK_PAC_FECV_03 => ("00000","00000","10000","11000","11110"),
  BLK_PAC_FECV_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_10 => ("00000","00001","00011","00111","00111"),
  BLK_PAC_FECV_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_14 => ("00000","10000","11000","11100","11100"),
  BLK_PAC_FECV_20 => ("01111","01111","01111","01111","01111"),
  BLK_PAC_FECV_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_22 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_24 => ("11110","11110","11110","11110","11110"),
  BLK_PAC_FECV_30 => ("00111","00111","00011","00001","00000"),
  BLK_PAC_FECV_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECV_34 => ("11100","11100","11000","10000","00000"),
  BLK_PAC_FECV_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECV_41 => ("01111","00011","00001","00000","00000"),
  BLK_PAC_FECV_42 => ("11111","11111","11111","00000","00000"),
  BLK_PAC_FECV_43 => ("11110","11000","10000","00000","00000"),
  BLK_PAC_FECV_44 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_00 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_01 => ("00000","00000","00011","00111","01111"),
  BLK_PAC_FECH_02 => ("00000","11111","11111","11111","11111"),
  BLK_PAC_FECH_03 => ("00000","00000","11000","11100","11110"),
  BLK_PAC_FECH_04 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_10 => ("00000","00001","00001","00011","00111"),
  BLK_PAC_FECH_11 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_12 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_13 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_14 => ("00000","10000","10000","11000","11100"),
  BLK_PAC_FECH_20 => ("00111","00111","00111","00111","00111"),
  BLK_PAC_FECH_21 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_22 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_23 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_24 => ("11100","11100","11100","11100","11100"),
  BLK_PAC_FECH_30 => ("00111","00011","00001","00001","00000"),
  BLK_PAC_FECH_31 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_32 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_33 => ("11111","11111","11111","11111","11111"),
  BLK_PAC_FECH_34 => ("11100","11000","10000","10000","00000"),
  BLK_PAC_FECH_40 => ("00000","00000","00000","00000","00000"),
  BLK_PAC_FECH_41 => ("01111","00111","00011","00000","00000"),
  BLK_PAC_FECH_42 => ("11111","11111","11111","11111","00000"),
  BLK_PAC_FECH_43 => ("11110","11100","11000","00000","00000"),
  BLK_PAC_FECH_44 => ("00000","00000","00000","00000","00000"),
  BLK_EYE_RED_CIM_00 => ("00001","10001","10001","11111","11111"),
  BLK_EYE_RED_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_CIM_02 => ("00010","00011","00011","11111","11111"),
  BLK_EYE_RED_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_RED_DIR_00 => ("01111","11111","11100","11100","11100"),
  BLK_EYE_RED_DIR_01 => ("00000","10001","00001","00001","00001"),
  BLK_EYE_RED_DIR_02 => ("11110","11111","11000","11000","11000"),
  BLK_EYE_RED_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_RED_BAI_00 => ("01111","11111","11111","11111","11000"),
  BLK_EYE_RED_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_BAI_02 => ("11110","11111","11111","11111","10001"),
  BLK_EYE_RED_BAI_10 => ("11000","01000","00000","00000","00000"),
  BLK_EYE_RED_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_BAI_12 => ("10001","10000","00000","00000","00000"),
  BLK_EYE_RED_ESQ_00 => ("01111","11111","00011","00011","00011"),
  BLK_EYE_RED_ESQ_01 => ("00000","10001","10000","10000","10000"),
  BLK_EYE_RED_ESQ_02 => ("11110","11111","00111","00111","00111"),
  BLK_EYE_RED_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_FAN_GRN_00 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_GRN_01 => ("00000","00111","01111","11111","11111"),
  BLK_FAN_GRN_02 => ("00000","11111","11111","11111","11111"),
  BLK_FAN_GRN_03 => ("00000","11000","11100","11110","11110"),
  BLK_FAN_GRN_04 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_GRN_10 => ("00001","00011","00011","00111","00111"),
  BLK_FAN_GRN_14 => ("00000","10000","10000","11000","11000"),
  BLK_FAN_GRN_20 => ("00111","00111","01111","01111","01111"),
  BLK_FAN_GRN_24 => ("11000","11000","11100","11100","11100"),
  BLK_FAN_GRN_30 => ("01111","01111","01111","01111","01111"),
  BLK_FAN_GRN_31 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_GRN_32 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_GRN_33 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_GRN_34 => ("11100","11100","11100","11100","11100"),
  BLK_FAN_GRN_40 => ("01111","01111","01111","00110","00000"),
  BLK_FAN_GRN_41 => ("10011","00001","00000","00000","00000"),
  BLK_FAN_GRN_42 => ("11111","11111","11110","01100","00000"),
  BLK_FAN_GRN_43 => ("10011","00001","00001","00000","00000"),
  BLK_FAN_GRN_44 => ("11100","11100","11100","11000","00000"),
  BLK_EYE_GRN_CIM_00 => ("10001","10001","10001","11111","11111"),
  BLK_EYE_GRN_CIM_01 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_02 => ("00011","00011","00011","11111","11111"),
  BLK_EYE_GRN_CIM_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_DIR_00 => ("11111","11111","11100","11100","11100"),
  BLK_EYE_GRN_DIR_01 => ("11111","11111","01111","01111","01111"),
  BLK_EYE_GRN_DIR_02 => ("11111","11111","11000","11000","11000"),
  BLK_EYE_GRN_DIR_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_DIR_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_DIR_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_BAI_00 => ("11111","11111","11111","11111","11000"),
  BLK_EYE_GRN_BAI_01 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_BAI_02 => ("11111","11111","11111","11111","10001"),
  BLK_EYE_GRN_BAI_10 => ("11000","11000","11111","11111","11111"),
  BLK_EYE_GRN_BAI_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_BAI_12 => ("10001","10001","11111","11111","11111"),
  BLK_EYE_GRN_ESQ_00 => ("11111","11111","00011","00011","00011"),
  BLK_EYE_GRN_ESQ_01 => ("11111","11111","11110","11110","11110"),
  BLK_EYE_GRN_ESQ_02 => ("11111","11111","00111","00111","00111"),
  BLK_EYE_GRN_ESQ_10 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_ESQ_11 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_GRN_ESQ_12 => ("11111","11111","11111","11111","11111"),
  BLK_EYE_BLK_CIM_00 => ("00001","10001","10001","11111","11111"),
  BLK_EYE_BLK_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_CIM_02 => ("00010","00011","00011","11111","11111"),
  BLK_EYE_BLK_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_DIR_00 => ("01111","11111","11100","11100","11100"),
  BLK_EYE_BLK_DIR_01 => ("00000","10001","00001","00001","00001"),
  BLK_EYE_BLK_DIR_02 => ("11110","11111","11000","11000","11000"),
  BLK_EYE_BLK_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_BAI_00 => ("01111","11111","11111","11111","11000"),
  BLK_EYE_BLK_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_BAI_02 => ("11110","11111","11111","11111","10001"),
  BLK_EYE_BLK_BAI_10 => ("11000","01000","00000","00000","00000"),
  BLK_EYE_BLK_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_BAI_12 => ("10001","10000","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_00 => ("01111","11111","00011","00011","00011"),
  BLK_EYE_BLK_ESQ_01 => ("00000","10001","10000","10000","10000"),
  BLK_EYE_BLK_ESQ_02 => ("11110","11111","00111","00111","00111"),
  BLK_EYE_BLK_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_FAN_VULN_00 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_01 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_02 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_03 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_04 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_10 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_11 => ("00000","00000","00000","00111","00111"),
  BLK_FAN_VULN_12 => ("00000","00000","00000","00001","00001"),
  BLK_FAN_VULN_13 => ("00000","00000","00000","11000","11000"),
  BLK_FAN_VULN_14 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_20 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_21 => ("00111","00000","00000","00000","00000"),
  BLK_FAN_VULN_22 => ("00001","00000","00000","00000","00000"),
  BLK_FAN_VULN_23 => ("11000","00000","00000","00000","00000"),
  BLK_FAN_VULN_24 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_30 => ("00000","00000","00011","00011","00000"),
  BLK_FAN_VULN_31 => ("11100","11100","00011","00011","00000"),
  BLK_FAN_VULN_32 => ("11110","11110","10011","10011","00000"),
  BLK_FAN_VULN_33 => ("01110","01110","10001","10001","00000"),
  BLK_FAN_VULN_34 => ("00000","00000","10000","10000","00000"),
  BLK_FAN_VULN_40 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_41 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_42 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_43 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_44 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_00 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_01 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_02 => ("00000","00000","00001","00011","00110"),
  BLK_MACA_03 => ("00000","00000","10000","00000","00000"),
  BLK_MACA_04 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_10 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_11 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_12 => ("00100","00000","00000","00000","00000"),
  BLK_MACA_13 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_14 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_20 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_21 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_22 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_23 => ("00000","00000","00000","00000","00110"),
  BLK_MACA_24 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_30 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_31 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_32 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_33 => ("00110","00100","00100","01000","00000"),
  BLK_MACA_34 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_40 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_41 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_42 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_43 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_44 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_00 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_01 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_02 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_03 => ("00000","00000","00011","00011","01111"),
  BLK_CEREJA_04 => ("00000","00000","10000","10000","10000"),
  BLK_CEREJA_10 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_11 => ("00000","00000","00000","00000","00001"),
  BLK_CEREJA_12 => ("00001","00110","01000","10000","00000"),
  BLK_CEREJA_13 => ("10001","00001","00010","00100","01000"),
  BLK_CEREJA_14 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_20 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_21 => ("00010","00000","00000","00000","00000"),
  BLK_CEREJA_22 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_23 => ("01000","01000","01000","00000","00000"),
  BLK_CEREJA_24 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_30 => ("00001","00000","00000","00000","00000"),
  BLK_CEREJA_31 => ("00000","10000","01000","00000","00000"),
  BLK_CEREJA_32 => ("00000","00000","00000","00010","00001"),
  BLK_CEREJA_33 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_34 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_40 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_41 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_42 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_43 => ("10000","00000","00000","00000","00000"),
  BLK_CEREJA_44 => ("00000","00000","00000","00000","00000"),
  OTHERS      => (OTHERS => (OTHERS => '0')));
  
  CONSTANT OVL_SPRITES_BLU: t_ovl_sprite5_vet := (
  BLK_EYE_GRN_CIM_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_CIM_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_GRN_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_GRN_DIR_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_GRN_DIR_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_DIR_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_GRN_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_GRN_BAI_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_GRN_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_BAI_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_GRN_BAI_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_BAI_12 => ("11111","11110","00000","00000","00000"),  
  BLK_EYE_GRN_ESQ_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_GRN_ESQ_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_GRN_ESQ_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_GRN_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_GRN_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_GRN_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_RED_CIM_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_RED_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_CIM_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_RED_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_RED_DIR_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_RED_DIR_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_DIR_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_RED_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_RED_BAI_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_RED_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_BAI_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_RED_BAI_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_BAI_12 => ("11111","11110","00000","00000","00000"),  
  BLK_EYE_RED_ESQ_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_RED_ESQ_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_RED_ESQ_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_RED_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_RED_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_RED_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_CIM_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_BLK_CIM_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_CIM_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_BLK_CIM_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_CIM_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_CIM_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_DIR_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_BLK_DIR_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_DIR_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_BLK_DIR_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_DIR_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_DIR_12 => ("11111","11110","00000","00000","00000"),
  BLK_EYE_BLK_BAI_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_BLK_BAI_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_BAI_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_BLK_BAI_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_BAI_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_BAI_12 => ("11111","11110","00000","00000","00000"),  
  BLK_EYE_BLK_ESQ_00 => ("01111","11111","11111","11111","11111"),
  BLK_EYE_BLK_ESQ_01 => ("00000","10001","10001","10001","10001"),
  BLK_EYE_BLK_ESQ_02 => ("11110","11111","11111","11111","11111"),
  BLK_EYE_BLK_ESQ_10 => ("11111","01111","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_11 => ("10001","00000","00000","00000","00000"),
  BLK_EYE_BLK_ESQ_12 => ("11111","11110","00000","00000","00000"),
  BLK_FAN_VULN_00 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_01 => ("00000","00111","01111","11111","11111"),
  BLK_FAN_VULN_02 => ("00000","11111","11111","11111","11111"),
  BLK_FAN_VULN_03 => ("00000","11000","11100","11110","11110"),
  BLK_FAN_VULN_04 => ("00000","00000","00000","00000","00000"),
  BLK_FAN_VULN_10 => ("00001","00011","00011","00111","00111"),
  BLK_FAN_VULN_11 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_12 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_13 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_14 => ("00000","10000","10000","11000","11000"),
  BLK_FAN_VULN_20 => ("00111","00111","01111","01111","01111"),
  BLK_FAN_VULN_21 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_22 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_23 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_24 => ("11000","11000","11100","11100","11100"),
  BLK_FAN_VULN_30 => ("01111","01111","01111","01111","01111"),
  BLK_FAN_VULN_31 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_32 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_33 => ("11111","11111","11111","11111","11111"),
  BLK_FAN_VULN_34 => ("11100","11100","11100","11100","11100"),
  BLK_FAN_VULN_40 => ("01111","01111","01111","00110","00000"),
  BLK_FAN_VULN_41 => ("10011","00001","00000","00000","00000"),
  BLK_FAN_VULN_42 => ("11111","11111","11110","01100","00000"),
  BLK_FAN_VULN_43 => ("10011","00001","00001","00000","00000"),
  BLK_FAN_VULN_44 => ("11100","11100","11100","11000","00000"),
  BLK_MACA_00 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_01 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_02 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_03 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_04 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_10 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_11 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_12 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_13 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_14 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_20 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_21 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_22 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_23 => ("00000","00000","00000","00000","00110"),
  BLK_MACA_24 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_30 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_31 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_32 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_33 => ("00110","00100","00100","01000","00000"),
  BLK_MACA_34 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_40 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_41 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_42 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_43 => ("00000","00000","00000","00000","00000"),
  BLK_MACA_44 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_00 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_01 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_02 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_03 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_04 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_10 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_11 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_12 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_13 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_14 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_20 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_21 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_22 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_23 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_24 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_30 => ("00001","00000","00000","00000","00000"),
  BLK_CEREJA_31 => ("00000","10000","01000","00000","00000"),
  BLK_CEREJA_32 => ("00000","00000","00000","00010","00001"),
  BLK_CEREJA_33 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_34 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_40 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_41 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_42 => ("00000","00000","00000","00000","00000"),
  BLK_CEREJA_43 => ("10000","00000","00000","00000","00000"),
  BLK_CEREJA_44 => ("00000","00000","00000","00000","00000"),
  OTHERS      => (OTHERS => (OTHERS => '0')));
END pac_sprites;
