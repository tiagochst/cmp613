LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.NUMERIC_STD.all;

ENTITY exemplo is
  PORT (    
    clk27M, reset_button      : in  STD_LOGIC;    
    red, green, blue          : out STD_LOGIC_vector(3 downto 0);
    hsync, vsync              : out STD_LOGIC);
END exemplo;

ARCHITECTURE comportamento of exemplo is
  SIGNAL rstn : STD_LOGIC;                      -- reset active low
                                        
  -- Interface com a mem�ria de v�deo do controlador
  SIGNAL we : STD_LOGIC;                        -- write enable ('1' p/ escrita)
  SIGNAL addr : integer range 0 to 12287;       -- ENDereco mem. vga
  SIGNAL pixel : STD_LOGIC_vector(2 downto 0);  -- valor de cor do pixel
  SIGNAL pixel_bit : STD_LOGIC;                 -- um bit do vetor acima

  -- Sinais dos contadores de linhas e colunas utilizados para percorrer
  -- as posi��es da mem�ria de v�deo (pixels) no momento de construir um quadro.
  SIGNAL line : integer range 0 to 95;          -- linha atual
  SIGNAL col : integer range 0 to 127;          -- coluna atual
  SIGNAL col_rstn : STD_LOGIC;                  -- reset do contador de colunas
  SIGNAL col_enable : STD_LOGIC;                -- enable do contador de colunas
  SIGNAL line_rstn : STD_LOGIC;                 -- reset do contador de linhas
  SIGNAL line_enable : STD_LOGIC;               -- enable do contador de linhas
  SIGNAL fim_escrita : STD_LOGIC;               -- '1' quando um quadro terminou de ser
                                                -- escrito na mem�ria de v�deo

  -- Especifica��o dos tipos e sinais da m�quina de estados de controle
  type estado_t is (show_splash, inicio, constroi_quadro, atualiza);
  SIGNAL estado: estado_t := show_splash;
  SIGNAL pr_estado: estado_t := show_splash;

  -- Sinais para um contador utilizado para atrasar a atualiza��o da
  -- posi��o da bola, a fim de evitar que a anima��o fique excessivamente
  -- veloz. Aqui utilizamos um contador de 0 a 270000, de modo que quando
  -- alimentado com um clock de 27MHz, ele demore 10ms para contar at� o final.
  SIGNAL contador : integer range 0 to 270000-1;
  SIGNAL timer : STD_LOGIC;                     -- vale '1' quando o contador chegar ao fim
  SIGNAL timer_rstn, timer_enable : STD_LOGIC;
  
  -- Defini��es de dados para o jogo
  subtype color3 is std_logic_vector(2 downto 0);
  type vcolor is array(0 to 3) of color3; 
  CONSTANT colors: vcolor :=                    -- cores de cada tipo de bloco tab_sym
  ("000", "001", "111", "100"); 
  
  type tab_sym is ('0', '1', '2', '3');         -- 0: vazio, 1; parede, 2: moeda, 3: porta
  type tab is array(0 to 95, 0 to 127) of tab_sym;
  
  --O cenario do jogo eh inicializado com todas as moedas e as paredes
  --As moedas v�o sendo removidas dessa estrutura de acordo com o jogo
  SIGNAL mapa:  tab := (
	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"01111111111111111111111111111111111111111000111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002002002002002002002001000100200200200200200200200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002001111111111002001111111111111002001000100200111111111111100200111111111100200100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01002001000000001002001000000000001002001000100200100000000000100200100000000100200100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01002001111111111002001111111111111002001111100200111111111111100200111111111100200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002002002002002002002002000200200200200200200200200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002001111111111002001111002001111111111111111111111100200111100200111111111100200100000000000000000000000000000000000000000000",
	"01000001000000001000001001000001000000000000000000000100000100100000100000000100000100000000000000000000000000000000000000000000",
	"01000001000000001000001001000001000000000000000000000100000100100000100000000100000100000000000000000000000000000000000000000000",
	"01002001111111111002001001002001111111111000111111111100200100100200111111111100200100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002001001002002002002001000100200200200200100100200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01111111111111111002001001111111111000001000100000111111111100100200111111111111111100000000000000000000000000000000000000000000",
	"00000000000000001000001000000000001000001000100000100000000000100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001000000000001000001000100000100000000000100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001111111111000001111100000111111111100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001000000000000000000000000000000000100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001000001111111110000011111111100000100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000013333310000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000010000010000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"01111111111111111002001111000001001111110000011111100100000111100200111111111111111100000000000000000000000000000000000000000000",
	"00000000000000000000000000000001001000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000001001000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000002000000000001001000000000000000100100000000000200000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000001001000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000001001000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000",
	"01111111111111111002001111000001001111111111111111100100000111100200111111111111111100000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000000000000000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000000000000000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001000001111111111111111111111100000100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001000000000000000000000000000000000100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000000000000000000000000000000000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001002001001000001111111111111111111111100000100100200100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000000000000000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"00000000000000001000001001000001000000000000000000000100000100100000100000000000000000000000000000000000000000000000000000000000",
	"01111111111111111002001111000001111111111000111111111100000111100200111111111111111100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002002002002002002002001000100200200200200200200200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000001000100000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002001111111111002001111111111111002001000100200111111111111100200111111111100200100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01000001000000001000001000000000001000001000100000100000000000100000100000000100000100000000000000000000000000000000000000000000",
	"01002001111111001002001111111111111002001111100200111111111111100200100111111100200100000000000000000000000000000000000000000000",
	"01000000000001001000000000000000000000000000000000000000000000000000100100000000000100000000000000000000000000000000000000000000",
	"01000000000001001000000000000000000000000000000000000000000000000000100100000000000100000000000000000000000000000000000000000000",
	"01002002002001001002002002002002002002000000000200200200200200200200100100200200200100000000000000000000000000000000000000000000",
	"01000000000001001000000000000000000000000000000000000000000000000000100100000000000100000000000000000000000000000000000000000000",
	"01000000000001001000000000000000000000000000000000000000000000000000100100000000000100000000000000000000000000000000000000000000",
	"01111111002001001002001111002001111111111111111111111100200111100200100100200111111100000000000000000000000000000000000000000000",
	"00000001000001001000001001000001000000000000000000000100000100100000100100000100000000000000000000000000000000000000000000000000",
	"00000001000001001000001001000001000000000000000000000100000100100000100100000100000000000000000000000000000000000000000000000000",
	"01111111002001111002001001002001111111111000111111111100200100100200111100200111111100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002001001002002002002001000100200200200200100100200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000001001000000000000001000100000000000000100100000000000000000000100000000000000000000000000000000000000000000",
	"01002001111111111111111001111111111002001000100200111111111100111111111111111100200100000000000000000000000000000000000000000000",
	"01000001000000000000000000000000001000001000100000100000000000000000000000000100000100000000000000000000000000000000000000000000",
	"01000001000000000000000000000000001000001000100000100000000000000000000000000100000100000000000000000000000000000000000000000000",
	"01002001111111111111111111111111111002001111100200111111111111111111111111111100200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01002002002002002002002002002002002002002000200200200200200200200200200200200200200100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"01111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
	);


BEGIN
  -- Controlador VGA (resolu��o 128 colunas por 96 linhas)
  -- Sinais:(aspect ratio 4:3). Os sinais que iremos utilizar para comunicar
  -- - write_clk (nosso clock)
  -- - write_enable ('1' quando queremos escrever um pixel)
  -- - write_addr (ENDere�o do pixel a escrever)
  -- - data_in (brilho do pixel RGB, 1 bit pra cada componente de cor)
  vga_controller: entity work.vgacon port map (
    clk27M       => clk27M,
    rstn         => '1',
    red          => red,
    green        => green,
    blue         => blue,
    hsync        => hsync,
    vsync        => vsync,
    write_clk    => clk27M,
    write_enable => we,
    write_addr   => addr,
    data_in      => pixel);

  -----------------------------------------------------------------------------
  -- Processos de varredura da tela
  -----------------------------------------------------------------------------
  
  -- purpose: Este processo conta o n�mero da coluna atual, quando habilitado
  --          pelo sinal "col_enable".
  -- type   : sequential
  -- inputs : clk27M, col_rstn
  -- outputs: col
  conta_coluna: PROCESS (clk27M, col_rstn)
  BEGIN  -- PROCESS conta_coluna
    IF col_rstn = '0' THEN                  -- asynchronous reset (active low)
      col <= 0;
    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
      IF col_enable = '1' THEN
        IF col = 127 THEN               -- conta de 0 a 127 (128 colunas)
          col <= 0;
        ELSE
          col <= col + 1;  
        END IF;
      END IF;
    END IF;
  END PROCESS conta_coluna;
    
  -- purpose: Este PROCESSo conta o n�mero da linha atual, quando habilitado
  --          pelo sinal "line_enable".
  -- type   : sequential
  -- inputs : clk27M, line_rstn
  -- outputs: line
  conta_linha: PROCESS (clk27M, line_rstn)
  BEGIN  -- PROCESS conta_linha
    IF line_rstn = '0' THEN                  -- asynchronous reset (active low)
      line <= 0;
    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
      -- o contador de linha s� incrementa quando o contador de colunas
      -- chegou ao fim (valor 127)
      IF line_enable = '1' and col = 127 THEN
        IF line = 95 THEN               -- conta de 0 a 95 (96 linhas)
          line <= 0;
        ELSE
          line <= line + 1;  
        END IF;        
      END IF;
    END IF;
  END PROCESS conta_linha;

  -- Este sinal � �til para informar nossa l�gica de controle quando
  -- o quadro terminou de ser escrito na mem�ria de v�deo, para que
  -- possamos avan�ar para o pr�ximo estado.
  fim_escrita <= '1' when (line = 95) and (col = 127)
                 ELSE '0'; 

  -----------------------------------------------------------------------------
  -- Abaixo est�o PROCESSos relacionados com a atualiza��o da posi��o da
  -- bola. Todos s�o controlados por sinais de enable de modo que a posi��o
  -- s� � de fato atualizada quando o controle (uma m�quina de estados)
  -- solicitar.
  -----------------------------------------------------------------------------

  -- purpose: Este PROCESSo ir� atualizar a coluna atual da bola,
  --          alterando sua posi��o no pr�ximo quadro a ser desenhado.
  -- type   : sequential
  -- inputs : clk27M, rstn
  -- outputs: pos_x
--  p_atualiza_pos_x: PROCESS (clk27M, rstn)
--    type direcao_t is (direita, esquerda);
--    VARIABLE direcao : direcao_t := direita;
--  BEGIN  -- PROCESS p_atualiza_pos_x
--    IF rstn = '0' THEN                  -- asynchronous reset (active low)
--      pos_x <= 0;
--    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
--      IF atualiza_pos_x = '1' THEN
--        IF direcao = direita THEN         
--          IF pos_x = 127 THEN
--            direcao := esquerda;  
--          ELSE
--            pos_x <= pos_x + 1;
--          END IF;        
--        ELSE  -- se a direcao � esquerda
--          IF pos_x = 0 THEN
--            direcao := direita;
--          ELSE
--            pos_x <= pos_x - 1;
--          END IF;
--        END IF;
--      END IF;
--    END IF;
--  END PROCESS p_atualiza_pos_x;
--
--  -- purpose: Este PROCESSo ir� atualizar a linha atual da bola,
--  --          alterando sua posi��o no pr�ximo quadro a ser desenhado.
--  -- type   : sequential
--  -- inputs : clk27M, rstn
--  -- outputs: pos_y
--  p_atualiza_pos_y: PROCESS (clk27M, rstn)
--    type direcao_t is (desce, sobe);
--    VARIABLE direcao : direcao_t := desce;
--  BEGIN  -- PROCESS p_atualiza_pos_x
--    IF rstn = '0' THEN                  -- asynchronous reset (active low)
--      pos_y <= 0;
--    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
--      IF atualiza_pos_y = '1' THEN
--        IF direcao = desce THEN         
--          IF pos_y = 95 THEN
--            direcao := sobe;  
--          ELSE
--            pos_y <= pos_y + 1;
--          END IF;        
--        ELSE  -- se a direcao � para subir
--          IF pos_y = 0 THEN
--            direcao := desce;
--          ELSE
--            pos_y <= pos_y - 1;
--          END IF;
--        END IF;
--      END IF;
--    END IF;
--  END PROCESS p_atualiza_pos_y;

  -----------------------------------------------------------------------------
  -- Brilho do pixel
  -----------------------------------------------------------------------------

  pixel_bit <= '1';
  pixel <= colors(0) WHEN mapa(line,col) = '0'
  ELSE     colors(1) WHEN mapa(line,col) = '1'
  ELSE     colors(2) WHEN mapa(line,col) = '2'
  ELSE     colors(3) WHEN mapa(line,col) = '3';
  
  -- O ENDere�o de mem�ria pode ser constru�do com essa f�rmula simples,
  -- a partir da linha e coluna atual
  addr  <= col + (128 * line);

  -----------------------------------------------------------------------------
  -- Processos que definem a FSM (finite state machine), nossa m�quina
  -- de estados de controle.
  -----------------------------------------------------------------------------

  -- purpose: Esta � a l�gica combinacional que calcula sinais de sa�da a partir
  --          do estado atual e alguns sinais de entrada (M�quina de Mealy).
  -- type   : combinational
  -- inputs : estado, fim_escrita, timer
  -- outputs: pr_estado, atualiza_pos_x, atualiza_pos_y, line_rstn,
  --          line_enable, col_rstn, col_enable, we, timer_enable, timer_rstn
  logica_mealy: PROCESS (estado, fim_escrita, timer)
  BEGIN  -- PROCESS logica_mealy
    case estado is
      when inicio         => IF timer = '1' THEN              
                               pr_estado <= constroi_quadro;
                             ELSE
                               pr_estado <= inicio;
                             END IF;
                             line_rstn      <= '0';  -- reset � active low!
                             line_enable    <= '0';
                             col_rstn       <= '0';  -- reset � active low!
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '1';  -- reset � active low!
                             timer_enable   <= '1';

      when constroi_quadro=> IF fim_escrita = '1' THEN
                               pr_estado <= atualiza;
                             ELSE
                               pr_estado <= constroi_quadro;
                             END IF;
                             line_rstn      <= '1';
                             line_enable    <= '1';
                             col_rstn       <= '1';
                             col_enable     <= '1';
                             we             <= '1';
                             timer_rstn     <= '0'; 
                             timer_enable   <= '0';

      when atualiza       => pr_estado <= inicio;
                             line_rstn      <= '1';
                             line_enable    <= '0';
                             col_rstn       <= '1';
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '0'; 
                             timer_enable   <= '0';

      when others         => pr_estado <= inicio;
                             line_rstn      <= '1';
                             line_enable    <= '0';
                             col_rstn       <= '1';
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '1'; 
                             timer_enable   <= '0';
      
    END case;
  END PROCESS logica_mealy;
  
  -- purpose: Avan�a a FSM para o pr�ximo estado
  -- type   : sequential
  -- inputs : clk27M, rstn, pr_estado
  -- outputs: estado
  seq_fsm: PROCESS (clk27M, rstn)
  BEGIN  -- PROCESS seq_fsm
    IF rstn = '0' THEN                  -- asynchronous reset (active low)
      estado <= inicio;
    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
      estado <= pr_estado;
    END IF;
  END PROCESS seq_fsm;

  -----------------------------------------------------------------------------
  -- Processos do contador utilizado para atrasar a anima��o (evitar
  -- que a atualiza��o de quadros fique excessivamente veloz).
  -----------------------------------------------------------------------------
  -- purpose: Incrementa o contador a cada ciclo de clock
  -- type   : sequential
  -- inputs : clk27M, timer_rstn
  -- outputs: contador, timer
  p_contador: PROCESS (clk27M, timer_rstn)
  BEGIN  -- PROCESS p_contador
    IF timer_rstn = '0' THEN            -- asynchronous reset (active low)
      contador <= 0;
    elsif clk27M'event and clk27M = '1' THEN  -- rising clock edge
      IF timer_enable = '1' THEN       
        IF contador = 270000 - 1 THEN
          contador <= 0;
        ELSE
          contador <=  contador + 1;        
        END IF;
      END IF;
    END IF;
  END PROCESS p_contador;

  -- purpose: Calcula o sinal "timer" que indica quando o contador chegou ao
  --          final
  -- type   : combinational
  -- inputs : contador
  -- outputs: timer
  p_timer: PROCESS (contador)
  BEGIN  -- PROCESS p_timer
    IF contador = 270000 - 1 THEN
      timer <= '1';
    ELSE
      timer <= '0';
    END IF;
  END PROCESS p_timer;

  -----------------------------------------------------------------------------
  -- Processos que sincronizam sinais ass�ncronos, de prefer�ncia com mais
  -- de 1 flipflop, para evitar metaestabilidade.
  -----------------------------------------------------------------------------
  
  -- purpose: Aqui sincronizamos nosso sinal de reset vindo do bot�o da DE1
  -- type   : sequential
  -- inputs : clk27M
  -- outputs: rstn
  build_rstn: PROCESS (clk27M)
    VARIABLE temp : STD_LOGIC;          -- flipflop intermediario
  BEGIN  -- PROCESS build_rstn
    IF clk27M'event and clk27M = '1' THEN  -- rising clock edge
      rstn <= temp;
      temp := reset_button;      
    END IF;
  END PROCESS build_rstn;

END comportamento;
