LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.PAC_DEFS.all;

ENTITY mem_mapa IS
	PORT 
	(
		clk		: IN STD_LOGIC;
		y_cor	: IN INTEGER range 0 to SCR_HGT - 1;
		x_cor	: IN INTEGER range 0 to SCR_WDT - 1;
		data	: IN tab_sym;
		we		: IN STD_LOGIC := '1';
		q		: OUT tab_sym;
		ledd : OUT STD_LOGIC
	);
END mem_mapa;

ARCHITECTURE rtl OF mem_mapa IS
	-- Build a 2-D array type FOR the RAM
	CONSTANT DATA_WIDTH: INTEGER := 4;
	type encoding_array is array(tab_sym) of std_logic_vector(DATA_WIDTH-1 downto 0);
	constant encode : encoding_array := ("0000", "0001", "0010", "0011", "0100");
	
	subtype word_t is std_logic_vector((DATA_WIDTH-1) downto 0);
	TYPE memory_t is array(SCR_HGT*SCR_WDT-1 downto 0) of word_t;
	
--	function init_ram
--		return memory_t is 
--		variable tmp : memory_t := (others => (others => '0'));
--	begin 
--		tmp := 		return tmp;
--	end init_ram;	 

	-- Declare the RAM SIGNAL and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	SIGNAL ram : memory_t := ("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0010","0100","0100","0100","0100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0010","0010","0010","0010","0010","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0001","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0001","0001","0011","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
		"0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000");
	attribute ram_init_file : string;
	attribute ram_init_file of ram : signal is "pacman.mif";

	-- Register to hold the address for (y,x) coordinates
	SIGNAL addr_reg, addr : INTEGER range 0 to SCR_HGT*SCR_WDT-1;

BEGIN
	PROCESS(clk, y_cor, x_cor)
	BEGIN
		addr <= y_cor*SCR_WDT + x_cor;
		
		IF(rising_edge(clk)) THEN
			IF(we = '1') THEN
				ram(addr) <= encode(data);
			END IF;

			-- Register the address FOR reading
			addr_reg <= addr;
		END IF;
	END PROCESS;

	--q <= ram(addr_reg);
	q <= ' ';
	
	ledd <= '1' WHEN ram(260) /= "0000"
	ELSE '0';
END rtl;
