LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY ram_64B IS
	PORT
	(
		clk       :IN STD_LOGIC ; 
		input     : IN STD_LOGIC_VECTOR (7 DOWNTO 0);  -- dados entrada
		output    : OUT STD_LOGIC_VECTOR (7 DOWNTO 0); -- saida
		address   : IN STD_LOGIC_VECTOR (5 DOWNTO 0);  -- endereco
		wren      : IN STD_LOGIC;                      -- W write-enable
		chipen    : IN STD_LOGIC;                      -- E chip-enable
		rden      : IN STD_LOGIC                       -- G read-enable
	);
END ram_64B;

ARCHITECTURE behav OF ram_64B IS
	SIGNAL address_sig : STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL clock_sig : STD_LOGIC ;
	SIGNAL clken_sig : STD_LOGIC ;
	SIGNAL data_sig: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL wren_sig,rden_sig: STD_LOGIC;
	SIGNAL q_sig : STD_LOGIC_VECTOR (7 DOWNTO 0);

COMPONENT ram1p IS
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		wren		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END COMPONENT ram1p;

BEGIN
	PROCESS(clk,wren,rden,chipen)
	 BEGIN
			IF(chipen = '1') THEN
				--write
				IF(wren='1' and rden ='0') THEN
					wren_sig <= '1';
					rden_sig <= '0';
				--read
				ELSIF(wren='0' and rden ='1') THEN
					wren_sig <= '0';
					rden_sig <= '1';
				--write and read -> nao 
				ELSE
					wren_sig <= '0';
					rden_sig <= '0';
				END IF;
			ELSE
				wren_sig <= '0';
				rden_sig <= '0';
			END IF;
	END PROCESS;

	PROCESS(q_sig, chipen, rden_sig) BEGIN
		IF(chipen = '1' and rden_sig = '1') THEN
			output<=q_sig;
		ELSE
			output<= (others=>'0');
		END IF;
	END PROCESS;

	ramp : ram1p PORT MAP (
			address,clk,input,wren_sig,q_sig
		);
END behav;