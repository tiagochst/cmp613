library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity alfa_char is 
port( code: IN STD_LOGIC_VECTOR(15 downto 0);
      alfa_code: OUT STD_LOGIC_VECTOR(6 downto 0));
end entity alfa_char;

architecture rtl of alfa_char is
begin
   process(code)
      begin
-- All choice expressions in a VHDL case statement must be constant
-- and unique.	Also, the case statement must be complete, or it must
-- include an others clause. 
      case (code) is
	  -- Sequential Statement(s)
	    when x"001c" =>
		  alfa_code <= "0001000"; --A
	    when x"0032" =>
		  alfa_code <= "0000011"; --B
	    when x"0021" =>
		  alfa_code <= "1000110"; --C
	    when x"0023" =>
		  alfa_code <= "0100001"; --D
	    when x"0024" =>
		  alfa_code <= "0000110"; --E
	    when x"002b" =>
		  alfa_code <= "0001110"; --F
	    when x"0034" =>
		  alfa_code <= "1000010"; --G
	    when x"0033" =>
		  alfa_code <= "0001011"; --h
	    when x"0043" =>
		  alfa_code <= "1001111"; --I
	    when x"003b" =>
		  alfa_code <= "1100000"; --J
	    when x"0042" =>
		  alfa_code <= "0001001"; --K
	    when x"004b" =>
		  alfa_code <= "1000111"; --L
	    when x"003a" =>
		  alfa_code <= "0000110"; --M
	    when x"0031" =>
		  alfa_code <= "0001110"; --N
	    when x"0044" =>
		  alfa_code <= "1000000"; --O
	    when x"004d" =>
		  alfa_code <= "0001100"; --P
	    when x"0015" =>
		  alfa_code <= "0011000"; --Q
	    when x"002d" =>
		  alfa_code <= "0101011"; --R
	    when x"001b" =>
		  alfa_code <= "0010010"; --S
	    when x"002c" =>
		  alfa_code <= "0001111"; --T
	    when x"003c" =>
		  alfa_code <= "1000001"; --U
	    when x"002a" =>
		  alfa_code <= "1100011"; --V
	    when x"001d" =>
		  alfa_code <= "0110000"; --W
	    when x"0022" =>
		  alfa_code <= "0001001"; --X
	    when x"0035" =>
		  alfa_code <= "0011001"; --Y
	    when x"001a" =>
		  alfa_code <= "0100100"; --Z
	    when x"0045" =>
		  alfa_code <= "1000000";
	    when x"0016" =>
		  alfa_code <= "1111001";
	    when x"001e" =>
		  alfa_code <= "0100100";
	    when x"0026" =>
		  alfa_code <= "0110000";
	    when x"0025" =>
		  alfa_code <= "0011001";
	    when x"002e" =>
		  alfa_code <= "0010010";
	    when x"0036" =>
		  alfa_code <= "0000010";
	    when x"003d" =>
		  alfa_code <= "1111000";
	    when x"003e" =>
		  alfa_code <= "0000000";
	    when x"0046" =>
		  alfa_code <= "0011000";
	    when others =>
		  alfa_code <="1111111";
      end case;
  end process;
END rtl;