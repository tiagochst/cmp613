LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.PAC_DEFS.all;

ENTITY mem_mapa IS
	PORT 
	(
		clk		: IN STD_LOGIC;
		y_cor	: IN INTEGER range 0 to SCR_HGT - 1;
		x_cor	: IN INTEGER range 0 to SCR_WDT - 1;
		data	: IN tab_sym;
		we		: IN STD_LOGIC := '1';
		q		: OUT tab_sym
	);
END mem_mapa;

ARCHITECTURE rtl OF mem_mapa IS
	-- Build a 2-D array type FOR the RAM
	TYPE memory_t is array(SCR_HGT*SCR_WDT-1 downto 0) of tab_sym;

	FUNCTION init_ram
		RETURN memory_t is 
		variable tmp : memory_t := (others =>' ');
	BEGIN 
		--O cen�rio do jogo � inicializado com todas as moedas e as paredes
		--As moedas v�o sendo removidas dessa estrutura de acordo com o jogo
		--O pacman e os fantasmas s�o desenhados separadamente sob essa tela
		tmp := (
	"                                                                                                                                "&
	"                                                                                                                                "&
	" 1111111111111111111111111111111111111111   1111111111111111111111111111111111111111                                            "&
	" 1                                      1   1                                      1                                            "&
	" 1                                      1   1                                      1                                            "& 
	" 1  2..2..2..2..2..2..2..2..2..2..2..2  1   1  2..2..2..2..2..2..2..2..2..2..2..2  1                                            "&
	" 1  .              .                 .  1   1  .                 .              .  1                                            "& 
	" 1  .              .                 .  1   1  .                 .              .  1                                            "&
	" 1  2  1111111111  2  1111111111111  2  1   1  2  1111111111111  2  1111111111  2  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  2  1        1  2  1           1  2  1   1  2  1           1  2  1        1  2  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  2  1111111111  2  1111111111111  2  11111  2  1111111111111  2  1111111111  2  1                                            "& 
	" 1  .              .                 .         .                 .              .  1                                            "& 
	" 1  .              .                 .         .                 .              .  1                                            "& 
	" 1  2..2..2..2..2..2..2..2..2..2..2..2..2...2..2..2..2..2..2..2..2..2..2..2..2..2  1                                            "& 
	" 1  .              .        .                           .        .              .  1                                            "& 
	" 1  .              .        .                           .        .              .  1                                            "& 
	" 1  2  1111111111  2  1111  2  11111111111111111111111  2  1111  2  1111111111  2  1                                            "& 
	" 1  .  1        1  .  1  1  .  1                     1  .  1  1  .  1        1  .  1                                            "& 
	" 1  .  1        1  .  1  1  .  1                     1  .  1  1  .  1        1  .  1                                            "& 
	" 1  2  1111111111  2  1  1  2  1111111111   1111111111  2  1  1  2  1111111111  2  1                                            "& 
	" 1  .              .  1  1  .           1   1           .  1  1  .              .  1                                            "& 
	" 1  .              .  1  1  .           1   1           .  1  1  .              .  1                                            "& 
	" 1  2..2..2..2..2..2  1  1  2..2..2..2  1   1  2..2..2..2  1  1  2..2..2..2..2..2  1                                            "& 
	" 1                 .  1  1           .  1   1  .           1  1  .                 1                                            "& 
	" 1                 .  1  1           .  1   1  .           1  1  .                 1                                            "& 
	" 1111111111111111  2  1  1111111111  .  1   1  .  1111111111  1  2  1111111111111111                                            "& 
	"                1  .  1           1  .  1   1  .  1           1  .  1                                                           "& 
	"                1  .  1           1  .  1   1  .  1           1  .  1                                                           "& 
	"                1  2  1  1111111111  .  11111  .  1111111111  1  2  1                                                           "& 
	"                1  .  1  1           .         .           1  1  .  1                                                           "& 
	"                1  .  1  1           .         .           1  1  .  1                                                           "& 
	"                1  2  1  1  .............................  1  1  2  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  2  1  1  .  111111111     111111111  .  1  1  2  1                                                           "& 
	"                1  .  1  1  .  1       1333331       1  .  1  1  .  1                                                           "& 
	"                1  .  1  1  .  1       1     1       1  .  1  1  .  1                                                           "& 
	" 1111111111111111  2  1111  .  1  111111     111111  1  .  1111  2  1111111111111111                                            "& 
	"                   .        .  1  1               1  1  .        .                                                              "& 
	"                   .        .  1  1               1  1  .        .                                                              "& 
	" ..................2.........  1  1               1  1  .........2..................                                            "& 
	"                   .        .  1  1               1  1  .        .                                                              "& 
	"                   .        .  1  1               1  1  .        .                                                              "& 
	" 1111111111111111  2  1111  .  1  11111111111111111  1  .  1111  2  1111111111111111                                            "& 
	"                1  .  1  1  .  1                     1  .  1  1  .  1                                                           "& 
	"                1  .  1  1  .  1                     1  .  1  1  .  1                                                           "& 
	"                1  2  1  1  .  11111111111111111111111  .  1  1  2  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  2  1  1  .............................  1  1  2  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  .  1  1  .                           .  1  1  .  1                                                           "& 
	"                1  2  1  1  .  11111111111111111111111  .  1  1  2  1                                                           "& 
	"                1  .  1  1  .  1                     1  .  1  1  .  1                                                           "& 
	"                1  .  1  1  .  1                     1  .  1  1  .  1                                                           "& 
	" 1111111111111111  2  1111  .  1111111111   1111111111  .  1111  2  1111111111111111                                            "& 
	" 1                 .        .           1   1           .        .                 1                                            "& 
	" 1                 .        .           1   1           .        .                 1                                            "& 
	" 1  2..2..2..2..2..2..2..2..2..2..2..2  1   1  2..2..2..2..2..2..2..2..2..2..2..2  1                                            "& 
	" 1  .              .                 .  1   1  .                 .              .  1                                            "& 
	" 1  .              .                 .  1   1  .                 .              .  1                                            "& 
	" 1  2  1111111111  2  1111111111111  2  1   1  2  1111111111111  2  1111111111  2  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  .  1        1  .  1           1  .  1   1  .  1           1  .  1        1  .  1                                            "& 
	" 1  2  1111111  1  2  1111111111111  2  11111  2  1111111111111  2  1  1111111  2  1                                            "& 
	" 1  .        1  1  .                 .         .                 .  1  1        .  1                                            "& 
	" 1  .        1  1  .                 .         .                 .  1  1        .  1                                            "& 
	" 1  2..2..2  1  1  2..2..2..2..2..2..2.........2..2..2..2..2..2..2  1  1  2..2..2  1                                            "& 
	" 1        .  1  1  .        .                           .        .  1  1  .        1                                            "& 
	" 1        .  1  1  .        .                           .        .  1  1  .        1                                            "& 
	" 1111111  2  1  1  2  1111  2  11111111111111111111111  2  1111  2  1  1  2  1111111                                            "& 
	"       1  .  1  1  .  1  1  .  1                     1  .  1  1  .  1  1  .  1                                                  "& 
	"       1  .  1  1  .  1  1  .  1                     1  .  1  1  .  1  1  .  1                                                  "& 
	" 1111111  2  1111  2  1  1  2  1111111111   1111111111  2  1  1  2  1111  2  1111111                                            "& 
	" 1        .        .  1  1  .           1   1           .  1  1  .        .        1                                            "& 
	" 1        .        .  1  1  .           1   1           .  1  1  .        .        1                                            "& 
	" 1  2..2..2..2..2..2  1  1  2..2..2..2  1   1  2..2..2..2  1  1  2..2..2..2..2..2  1                                            "& 
	" 1  .                 1  1           .  1   1  .           1  1                 .  1                                            "& 
	" 1  .                 1  1           .  1   1  .           1  1                 .  1                                            "& 
	" 1  2  1111111111111111  1111111111  2  1   1  2  1111111111  1111111111111111  2  1                                            "& 
	" 1  .  1                          1  .  1   1  .  1                          1  .  1                                            "& 
	" 1  .  1                          1  .  1   1  .  1                          1  .  1                                            "& 
	" 1  2  1111111111111111111111111111  2  11111  2  1111111111111111111111111111  2  1                                            "& 
	" 1  .                                .         .                                .  1                                            "& 
	" 1  .                                .         .                                .  1                                            "& 
	" 1  2..2..2..2..2..2..2..2..2..2..2..2..2...2..2..2..2..2..2..2..2..2..2..2..2..2  1                                            "& 
	" 1                                                                                 1                                            "& 
	" 1                                                                                 1                                            "& 
	" 11111111111111111111111111111111111111111111111111111111111111111111111111111111111                                            "& 
	"                                                                                                                                "& 
	"                                                                                                                                "& 
	"                                                                                                                                "
	);
		RETURN tmp;
	END init_ram;	 

	-- Declare the RAM SIGNAL and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	SIGNAL ram : memory_t := init_ram;

	-- Register to hold the address for (y,x) coordinates
	SIGNAL addr_reg, addr : INTEGER range 0 to SCR_HGT*SCR_WDT-1;

BEGIN
	PROCESS(clk, y_cor, x_cor)
	BEGIN
		addr <= y_cor*SCR_WDT + x_cor;
		
		IF(rising_edge(clk)) THEN
			IF(we = '1') THEN
				ram(addr) <= data;
			END IF;

			-- Register the address FOR reading
			addr_reg <= addr;
		END IF;
	END PROCESS;

	q <= ram(addr_reg);
END rtl;
